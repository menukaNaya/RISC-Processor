// Define the stimulus module (no ports)
module stimulus;

	// Declare variables to be connected
	// to inputs
	reg IN0, IN1;
	reg S0;
	
	// Declare output wire
	wire OUTPUT;
	
	// Instantiate the multiplexer
	mux2_to_1 mymux(OUTPUT, IN0, IN1, S0);
	
	// Stimulate the inputs
	// Define the stimulus module (no ports)
	initial
	begin
		// set input lines
		IN0 = 1; IN1 = 0;
		#1 $display("IN0= %b, IN1= %b \n",IN0,IN1);
		// choose IN0
		S0 = 0;
		#1 $display("S0 = %b, OUTPUT = %b \n", S0, OUTPUT);
		// choose IN1
		S0 = 1;
		#1 $display("S0 = %b, OUTPUT = %b \n", S0, OUTPUT);
		
	end
	
endmodule


// Module 4-to-1 multiplexer. Port list is taken exactly from
// the I/O diagram.
module mux2_to_1 (out, i0, i1, s0);
	
	// Port declarations from the I/O diagram
	output out;
	input i0, i1;
	input s0;

	reg tempout;
	
	always @(s0,i0,i1)
	begin	
	
	if (s0==1'b0)
		tempout = i0;
	else
		tempout = i1;	
	end	
	
	assign out=tempout;
	
endmodule
